module main

import ui

fn btn_help_click(b voidptr) {
	ui.message_box('Built with V UI')
}